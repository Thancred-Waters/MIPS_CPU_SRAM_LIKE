`define CR_STATUS   5'b01100
`define CR_COMPARE  5'b01011
`define CR_CAUSE    5'b01101
`define CR_EPC      5'b01110
`define CR_COUNT    5'b01001
`define CR_BADVADDR 5'b01000

`define EX_INT  5'h00
`define EX_ADEL 5'h04
`define EX_ADES 5'h05
`define EX_OV   5'h0c
`define EX_SYS  5'h08
`define EX_BP   5'h09
`define EX_RI   5'h0a